module jb_control_unit (
    input  logic    stall_F,
    input  logic    R,
    input  logic    zero,
    output logic    stall_EX,
    output logic    pc_src
)



endmodule