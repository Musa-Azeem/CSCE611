module jb_control_unit (
    input logic     stall_F,
    output logic    stall_EX,

)
endmodule